library verilog;
use verilog.vl_types.all;
entity seq is
    generic(
        S_IF1           : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        \S_IF2\         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        \S_IMM1\        : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        \S_IMM2\        : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        \S_MR1\         : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        \S_MR2\         : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        \S_DISP\        : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        \S_IN\          : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        \S_IACK\        : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        \S_MW1\         : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi0);
        \S_MW2\         : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi1);
        \S_OUT\         : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1)
    );
    port(
        data_in         : in     vl_logic_vector(7 downto 0);
        busreq          : in     vl_logic;
        waitreq         : in     vl_logic;
        intreq          : in     vl_logic;
        nmireq          : in     vl_logic;
        reset_in        : in     vl_logic;
        clk             : in     vl_logic;
        intack_out      : out    vl_logic;
        nmiack_out      : out    vl_logic;
        busack_out      : out    vl_logic;
        iff2_out        : out    vl_logic;
        icb_out         : out    vl_logic;
        idd_out         : out    vl_logic;
        ied_out         : out    vl_logic;
        ifd_out         : out    vl_logic;
        inst_reg        : out    vl_logic_vector(7 downto 0);
        start           : out    vl_logic;
        mreq            : out    vl_logic;
        iorq            : out    vl_logic;
        rd              : out    vl_logic;
        wr              : out    vl_logic;
        imm1            : in     vl_logic;
        imm2            : in     vl_logic;
        mr1             : in     vl_logic;
        mr2             : in     vl_logic;
        mw1             : in     vl_logic;
        mw2             : in     vl_logic;
        disp            : in     vl_logic;
        i_in            : in     vl_logic;
        i_out           : in     vl_logic;
        i_eidi          : in     vl_logic;
        i_im            : in     vl_logic;
        retin           : in     vl_logic;
        i43             : in     vl_logic_vector(1 downto 0);
        g_if            : out    vl_logic;
        g_imm2          : out    vl_logic;
        g_mr1           : out    vl_logic;
        g_mr2           : out    vl_logic;
        g_mw1           : out    vl_logic;
        g_mw2           : out    vl_logic;
        g_disp          : out    vl_logic;
        g_in            : out    vl_logic;
        g_out           : out    vl_logic;
        g_iack          : out    vl_logic;
        sgate           : out    vl_logic;
        s_if            : out    vl_logic;
        s_if2           : out    vl_logic;
        s_imm1          : out    vl_logic;
        s_imm2          : out    vl_logic;
        s_mr1           : out    vl_logic;
        s_mr2           : out    vl_logic;
        s_mw1           : out    vl_logic;
        s_mw2           : out    vl_logic;
        s_disp          : out    vl_logic;
        s_in            : out    vl_logic;
        s_out           : out    vl_logic;
        s_iack          : out    vl_logic;
        m1              : out    vl_logic;
        intmode         : out    vl_logic_vector(1 downto 0);
        i_halt          : in     vl_logic;
        eschalt         : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of S_IF1 : constant is 1;
    attribute mti_svvh_generic_type of \S_IF2\ : constant is 1;
    attribute mti_svvh_generic_type of \S_IMM1\ : constant is 1;
    attribute mti_svvh_generic_type of \S_IMM2\ : constant is 1;
    attribute mti_svvh_generic_type of \S_MR1\ : constant is 1;
    attribute mti_svvh_generic_type of \S_MR2\ : constant is 1;
    attribute mti_svvh_generic_type of \S_DISP\ : constant is 1;
    attribute mti_svvh_generic_type of \S_IN\ : constant is 1;
    attribute mti_svvh_generic_type of \S_IACK\ : constant is 1;
    attribute mti_svvh_generic_type of \S_MW1\ : constant is 1;
    attribute mti_svvh_generic_type of \S_MW2\ : constant is 1;
    attribute mti_svvh_generic_type of \S_OUT\ : constant is 1;
end seq;
